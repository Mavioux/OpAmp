** Profile: "SCHEMATIC1-simulation"  [ F:\Users\Mavioux\Orcad Projects\telestikos enisxyths-pspicefiles\schematic1\simulation.sim ] 

** Creating circuit file "simulation.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../telestikos enisxyths-pspicefiles/telestikos enisxyths.lib" 
* From [PSPICE NETLIST] section of F:\CADENCE\WORKING DIRECTORY\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 4200us 0 SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
