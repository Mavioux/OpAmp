** Profile: "SCHEMATIC1-ac sweer"  [ F:\Users\Mavioux\Orcad Projects\telestikos enisxyths-pspicefiles\schematic1\ac sweer.sim ] 

** Creating circuit file "ac sweer.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../telestikos enisxyths-pspicefiles/telestikos enisxyths.lib" 
* From [PSPICE NETLIST] section of F:\CADENCE\WORKING DIRECTORY\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 0.1 10g
.TEMP 0 10 20 30 40 50 60
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
